module imem #(parameter N = 32)
				(input logic [5:0] addr,
				 output logic [N-1:0] q);
	// Here goes the implementation of imem
	// Ver tema de arreglos para almacenamiento de la info necesaria
endmodule